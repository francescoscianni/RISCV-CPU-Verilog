module alu (
    input [31:0] a,
    input [31:0] b,
    input [2:0] alucontrol,
    output reg [31:0] result,
    output zero
);

assign zero = (result == 32'd0);

always @(*) begin
    case (alucontrol)
        3'b000: result = a + b;   // ADD
        3'b001: result = a - b;   // SUB
        3'b010: result = a << b[4:0];   // SLL
        3'b011: result = a < b ? 32'd1:32'd0 ;   // SLT
        3'b100: result = a^b; //XOR
        3'b101: result = a >> b[4:0]; //SRL
        3'b110: result = a | b; //OR
        3'b111: result = a & b; //AND
    endcase
end

endmodule
//cpu.v alu.v cu.v mux2_1.v extend.v mux3_1.v ram.v regfile.v regnbit.v