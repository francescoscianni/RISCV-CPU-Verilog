module AND (
    input wire A,    // Input A
    input wire B,    // Input B
    output wire Y    // Out Y = A AND B
);
    assign Y = A & B; 
endmodule